----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:03:27 04/23/2012 
-- Design Name: 
-- Module Name:    SpriteGpu - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SpriteGpu is
    Port ( 	clk : in  STD_LOGIC;
				x : in  integer;
				y : in  integer;
				spriteVgaRed: out  std_logic_vector(2 downto 0);					
				spriteVgaGreen: out  std_logic_vector(2 downto 0);		
				spriteVgaBlue: out  std_logic_vector(2 downto 1);
				collision: out std_logic;
				spriteDetected: out std_logic;
				rst : in  STD_LOGIC;
				jump: in std_logic;
				duck: in std_logic;
				move_box: in std_logic;
				put_box: in std_logic;
				next_box: in std_logic;
				split_legs: in std_logic);
end SpriteGpu;


architecture Behavioral of SpriteGpu is

subtype elements is std_logic_vector(31 downto 0);
type bit_array is array (0 to 31) of elements;
type gubb_array is array (0 to 64) of elements;
subtype test is integer  range 0 to 800;
type position is array (0 to 7) of test;
signal sprite_brick : bit_array ;
signal sprite_gubbe:  gubb_array;
signal sprite_gubbe_aktiv:  gubb_array;
signal sprite_gubbe_jump:  gubb_array;
signal sprite_gubbe_duck:  gubb_array;
signal sprite_gubbe_split:  gubb_array;
signal x_pos : position;
signal y_pos : position;

signal spriteSize : integer := 32;
signal gubbSize : integer := 64;
signal btnuPressed: std_logic;
begin


sprite_brick( 0) <= "11111111111111111111111111111111"; 
sprite_brick( 1) <= "10010010010010000100100100100101"; 
sprite_brick( 2) <= "11001001001001001001001001001001"; 
sprite_brick( 3) <= "10100100100100100100100100100101";
sprite_brick( 4) <= "10010010010010000100100100100101"; 
sprite_brick( 5) <= "11001001001001001001001001001001"; 
sprite_brick( 6) <= "10100100100100100100100100100101"; 
sprite_brick( 7) <= "10010010010010000100100100100101"; 
sprite_brick( 8) <= "11001001001001001001001001001001"; 
sprite_brick( 9) <= "10100100100100100100100100100101"; 
sprite_brick(10) <= "10010010010010000100100100100101"; 
sprite_brick(11) <= "11001001001001001001001001001001"; 
sprite_brick(12) <= "10100100100100100100100100100101"; 
sprite_brick(13) <= "10010010010010000100100100100101"; 
sprite_brick(14) <= "11001001001001001001001001001001"; 
sprite_brick(15) <= "10100100100100100100100100100101";
sprite_brick(16) <= "10010010010010000100100100100101"; 
sprite_brick(17) <= "11001001001001001001001001001001"; 
sprite_brick(18) <= "10100100100100100100100100100101"; 
sprite_brick(19) <= "10010010010010000100100100100101"; 
sprite_brick(20) <= "11001001001001001001001001001001"; 
sprite_brick(21) <= "10100100100100100100100100100101"; 
sprite_brick(22) <= "10010010010010000100100100100101"; 
sprite_brick(23) <= "11001001001001001001001001001001"; 
sprite_brick(24) <= "10100100100100100100100100100101"; 
sprite_brick(25) <= "10010010010010000100100100100101"; 
sprite_brick(26) <= "11001001001001001001001001001001"; 
sprite_brick(27) <= "10100100100100100100100100100101"; 
sprite_brick(28) <= "10010010010010000100100100100101"; 
sprite_brick(29) <= "11001001001001001001001001001001"; 
sprite_brick(30) <= "10100100100100100100100100100101"; 
sprite_brick(31) <= "11111111111111111111111111111111";  

sprite_gubbe( 0) <= "00000111000111000000011100011100";
sprite_gubbe( 1) <= "00001100000011100000110000001110";
sprite_gubbe( 2) <= "00011001110001110000110000001110";
sprite_gubbe( 3) <= "00110011111001110000110000001110";
sprite_gubbe( 4) <= "00110011111001110000110000001110";
sprite_gubbe( 5) <= "01110011110001110000110000001110";
sprite_gubbe( 6) <= "01110001100011100000110000001110";
sprite_gubbe( 7) <= "01111111111111100000110000001110";
sprite_gubbe( 8) <= "01111111111111100000110000001110";
sprite_gubbe( 9) <= "01111111111111000000110000001110";
sprite_gubbe(10) <= "01111111111111000000110000001110";
sprite_gubbe(11) <= "00111111111111000000110000001110";
sprite_gubbe(12) <= "00111111111111000000110000001110";
sprite_gubbe(13) <= "00111111111111000000110000001110";
sprite_gubbe(14) <= "00011111111110000000110000001110";
sprite_gubbe(15) <= "00011111111110000000110000001110";
sprite_gubbe(16) <= "00011111111110000000110000001110";
sprite_gubbe(17) <= "00011111111110000000110000001110";
sprite_gubbe(18) <= "00011111111110000000110000001110";
sprite_gubbe(19) <= "00011111011111000000110000001110";
sprite_gubbe(20) <= "00111110001111100000110000001110";
sprite_gubbe(21) <= "00111110001111100000110000001110";
sprite_gubbe(22) <= "00111110001111100000110000001110";
sprite_gubbe(23) <= "00111110001111100000110000001110";
sprite_gubbe(24) <= "01111100001111100000110000001110";
sprite_gubbe(25) <= "11111000001111000000110000001110";
sprite_gubbe(26) <= "11111000001110000000110000001110";
sprite_gubbe(27) <= "11110000001110000000110000001110";
sprite_gubbe(28) <= "11110000001110000000110000001110";
sprite_gubbe(29) <= "11110000001111000000110000001110";
sprite_gubbe(30) <= "11111110001111110000110000001110";
sprite_gubbe(31) <= "11111110001111110000110000001110";
sprite_gubbe(32) <= "00000111000111000000011100011100";
sprite_gubbe(33) <= "00001100000011100000110000001110";
sprite_gubbe(34) <= "00011001110001110000110000001110";
sprite_gubbe(35) <= "00110011111001110000110000001110";
sprite_gubbe(36) <= "00110011111001110000110000001110";
sprite_gubbe(37) <= "01110011110001110000110000001110";
sprite_gubbe(38) <= "01110001100011100000110000001110";
sprite_gubbe(39) <= "01111111111111100000110000001110";
sprite_gubbe(40) <= "01111111111111100000110000001110";
sprite_gubbe(41) <= "01111111111111000000110000001110";
sprite_gubbe(42) <= "01111111111111000000110000001110";
sprite_gubbe(43) <= "00111111111111000000110000001110";
sprite_gubbe(44) <= "00111111111111000000110000001110";
sprite_gubbe(45) <= "00111111111111000000110000001110";
sprite_gubbe(46) <= "00011111111110000000110000001110";
sprite_gubbe(47) <= "00011111111110000000110000001110";
sprite_gubbe(48) <= "00011111111110000000110000001110";
sprite_gubbe(49) <= "00011111111110000000110000001110";
sprite_gubbe(50) <= "00011111111110000000110000001110";
sprite_gubbe(51) <= "00011111011111000000110000001110";
sprite_gubbe(52) <= "00111110001111100000110000001110";
sprite_gubbe(53) <= "00111110001111100000110000001110";
sprite_gubbe(54) <= "00111110001111100000110000001110";
sprite_gubbe(55) <= "00111110001111100000110000001110";
sprite_gubbe(56) <= "01111100001111100000110000001110";
sprite_gubbe(57) <= "11111000001111000000110000001110";
sprite_gubbe(58) <= "11111000001110000000110000001110";
sprite_gubbe(59) <= "11110000001110000000110000001110";
sprite_gubbe(60) <= "11110000001110000000110000001110";
sprite_gubbe(61) <= "11110000001111000000110000001110";
sprite_gubbe(62) <= "11111110001111110000110000001110";
sprite_gubbe(63) <= "11111110001111110000110000001110";

sprite_gubbe_jump( 0) <= "00000111000111000000011100011100";
sprite_gubbe_jump( 1) <= "00001100000011100000110000001110";
sprite_gubbe_jump( 2) <= "00011001110001110000110000001110";
sprite_gubbe_jump( 3) <= "00110011111001110000110000001110";
sprite_gubbe_jump( 4) <= "00110011111001110111111111111110";
sprite_gubbe_jump( 5) <= "01110011110001110000110000001110";
sprite_gubbe_jump( 6) <= "01110001100011100000110000001110";
sprite_gubbe_jump( 7) <= "01111111111111100000110000001110";
sprite_gubbe_jump( 8) <= "01111111111111100000110000001110";
sprite_gubbe_jump( 9) <= "01111111111111000000110000001110";
sprite_gubbe_jump(10) <= "01111111111111001111111111101110";
sprite_gubbe_jump(11) <= "00000000000000000000110000001110";
sprite_gubbe_jump(12) <= "00111111111111000000110000001110";
sprite_gubbe_jump(13) <= "00111111111111000000110000001110";
sprite_gubbe_jump(14) <= "00011111111110000000110000001110";
sprite_gubbe_jump(15) <= "00011111111110000000110000001110";
sprite_gubbe_jump(16) <= "00011111111110001111111100001110";
sprite_gubbe_jump(17) <= "00011111111110000000110000001110";
sprite_gubbe_jump(18) <= "00011111111110000000110000001110";
sprite_gubbe_jump(19) <= "00011111011111000000110000001110";
sprite_gubbe_jump(20) <= "00111110001111100000110000001110";
sprite_gubbe_jump(21) <= "00111110001111100000110000001110";
sprite_gubbe_jump(22) <= "00111111111111111111000000001110";
sprite_gubbe_jump(23) <= "00111110001111100000110000001110";
sprite_gubbe_jump(24) <= "01111100001111100000110000001110";
sprite_gubbe_jump(25) <= "11111111111111111111111111111110";
sprite_gubbe_jump(26) <= "11111000001110000000110000001110";
sprite_gubbe_jump(27) <= "11111111111111111111111111111110";
sprite_gubbe_jump(28) <= "11110000001110000000110000001110";
sprite_gubbe_jump(29) <= "11110000001111000000110000001110";
sprite_gubbe_jump(30) <= "11111110001111110000110000001110";
sprite_gubbe_jump(31) <= "11111110111111111111110000001110";
sprite_gubbe_jump(32) <= "00000111000111000000011100011100";
sprite_gubbe_jump(33) <= "00001100000011100000110000001110";
sprite_gubbe_jump(34) <= "00011001110001110000110000001110";
sprite_gubbe_jump(35) <= "00110011111001110000110000001110";
sprite_gubbe_jump(36) <= "00110011111001110000110000001110";
sprite_gubbe_jump(37) <= "01110011110001110000110000001110";
sprite_gubbe_jump(38) <= "01110001100011100000110000001110";
sprite_gubbe_jump(39) <= "01111111111111100000110000001110";
sprite_gubbe_jump(40) <= "01111111111111100000110000001110";
sprite_gubbe_jump(41) <= "01111111111111000000110000001110";
sprite_gubbe_jump(42) <= "01111111111111000000110000001110";
sprite_gubbe_jump(43) <= "00111111111111000000110000001110";
sprite_gubbe_jump(44) <= "00111111111111000000110000001110";
sprite_gubbe_jump(45) <= "00111111111111000000110000001110";
sprite_gubbe_jump(46) <= "00011111111110000000110000001110";
sprite_gubbe_jump(47) <= "00011111111110111111111111111110";
sprite_gubbe_jump(48) <= "00011111111110000000110000001110";
sprite_gubbe_jump(49) <= "00011111111110111111111111111110";
sprite_gubbe_jump(50) <= "00011100111111111111111111111110";
sprite_gubbe_jump(51) <= "00011111011111111111111100001110";
sprite_gubbe_jump(52) <= "00111110001111100000110000001110";
sprite_gubbe_jump(53) <= "00111110001111100000110000001110";
sprite_gubbe_jump(54) <= "00111110001111101111111111111110";
sprite_gubbe_jump(55) <= "00111110001111100000110000001110";
sprite_gubbe_jump(56) <= "01111100001111100000110000001110";
sprite_gubbe_jump(57) <= "11111000001111000000110000001110";
sprite_gubbe_jump(58) <= "11111000001110001111110000001110";
sprite_gubbe_jump(59) <= "11110000001110000000110000001110";
sprite_gubbe_jump(60) <= "11110000001110000000110000001110";
sprite_gubbe_jump(61) <= "11110000001111000000110000001110";
sprite_gubbe_jump(62) <= "11111110001111110000110000001110";
sprite_gubbe_jump(63) <= "11111110001111110000110000001110";

sprite_gubbe_duck( 0) <= "11110001110001111111000111000111";
sprite_gubbe_duck( 1) <= "11110011111100111110001111110010";
sprite_gubbe_duck( 2) <= "11000110011100011111001111110010";
sprite_gubbe_duck( 3) <= "11001100001110011111001111110010";
sprite_gubbe_duck( 4) <= "11001100001110010000000000000000";
sprite_gubbe_duck( 5) <= "00011100001100011111001111110010";
sprite_gubbe_duck( 6) <= "00011100011000111110001111110010";
sprite_gubbe_duck( 7) <= "00000000000000011110001111110010";
sprite_gubbe_duck( 8) <= "00000000000000011110001111110010";
sprite_gubbe_duck( 9) <= "00000000000001111111001111110010";
sprite_gubbe_duck(10) <= "00000000000001110000000000100010";
sprite_gubbe_duck(11) <= "11111111111111111111001111110010";
sprite_gubbe_duck(12) <= "11000000000000111111001111110010";
sprite_gubbe_duck(13) <= "11000000000000111111001111110010";
sprite_gubbe_duck(14) <= "11000000000001111110001111110010";
sprite_gubbe_duck(15) <= "11000000000001111110001111110010";
sprite_gubbe_duck(16) <= "11000000000001100000000011110010";
sprite_gubbe_duck(17) <= "11000000000001111110001111110010";
sprite_gubbe_duck(18) <= "11000000000001111110001111110010";
sprite_gubbe_duck(19) <= "11000001000001111111001111110010";
sprite_gubbe_duck(20) <= "11000011100000111110001111110010";
sprite_gubbe_duck(21) <= "11000011100000111110001111110010";
sprite_gubbe_duck(22) <= "11000000000000000000111111110010";
sprite_gubbe_duck(23) <= "11000011100000111110001111110010";
sprite_gubbe_duck(24) <= "00000111110000111110001111110010";
sprite_gubbe_duck(25) <= "00000000000000000000000000000010";
sprite_gubbe_duck(26) <= "00001111100011111110001111110010";
sprite_gubbe_duck(27) <= "00000000000000000000000000000010";
sprite_gubbe_duck(28) <= "00001111110011111110001111110010";
sprite_gubbe_duck(29) <= "00001111110000111111001111110010";
sprite_gubbe_duck(30) <= "00000011100000001111001111110010";
sprite_gubbe_duck(31) <= "00000010000000000000001111110010";
sprite_gubbe_duck(32) <= "00000000000000000000000000000000";
sprite_gubbe_duck(33) <= "00000000000000000000000000000000";
sprite_gubbe_duck(34) <= "00000000000000000000000000000000";
sprite_gubbe_duck(35) <= "00000000000000000000000000000000";
sprite_gubbe_duck(36) <= "00000000000000000000000000000000";
sprite_gubbe_duck(37) <= "00000000000000000000000000000000";
sprite_gubbe_duck(38) <= "00000000000000000000000000000000";
sprite_gubbe_duck(39) <= "00000000000000000000000000000000";
sprite_gubbe_duck(40) <= "00000000000000000000000000000000";
sprite_gubbe_duck(41) <= "00000000000000000000000000000000";
sprite_gubbe_duck(42) <= "00000000000000000000000000000000";
sprite_gubbe_duck(43) <= "00000000000000000000000000000000";
sprite_gubbe_duck(44) <= "00000000000000000000000000000000";
sprite_gubbe_duck(45) <= "00000000000000000000000000000000";
sprite_gubbe_duck(46) <= "00000000000000000000000000000000";
sprite_gubbe_duck(47) <= "00000000000000000000000000000000";
sprite_gubbe_duck(48) <= "00000000000000000000000000000000";
sprite_gubbe_duck(49) <= "00000000000000000000000000000000";
sprite_gubbe_duck(50) <= "00000000000000000000000000000000";
sprite_gubbe_duck(51) <= "00000000000000000000000000000000";
sprite_gubbe_duck(52) <= "00000000000000000000000000000000";
sprite_gubbe_duck(53) <= "00000000000000000000000000000000";
sprite_gubbe_duck(54) <= "00000000000000000000000000000000";
sprite_gubbe_duck(55) <= "00000000000000000000000000000000";
sprite_gubbe_duck(56) <= "00000000000000000000000000000000";
sprite_gubbe_duck(57) <= "00000000000000000000000000000000";
sprite_gubbe_duck(58) <= "00000000000000000000000000000000";
sprite_gubbe_duck(59) <= "00000000000000000000000000000000";
sprite_gubbe_duck(60) <= "00000000000000000000000000000000";
sprite_gubbe_duck(61) <= "00000000000000000000000000000000";
sprite_gubbe_duck(62) <= "00000000000000000000000000000000";
sprite_gubbe_duck(63) <= "00000000000000000000000000000000";

sprite_gubbe_split( 0) <= "11111111111111111111111111111111";
sprite_gubbe_split( 1) <= "11110011111100111111111111110010";
sprite_gubbe_split( 2) <= "11111110011111111111001111110010";
sprite_gubbe_split( 3) <= "11001111101110011111001111110010";
sprite_gubbe_split( 4) <= "11001111101110011111111111111110";
sprite_gubbe_split( 5) <= "11111111101111111111001111110010";
sprite_gubbe_split( 6) <= "11111111111111111111111111110010";
sprite_gubbe_split( 7) <= "11111111111111111111111111110010";
sprite_gubbe_split( 8) <= "11111111111111111111111111110010";
sprite_gubbe_split( 9) <= "11111111111101111111001111110010";
sprite_gubbe_split(10) <= "11111111111101111111111110111110";
sprite_gubbe_split(11) <= "11111111111111111111001111110010";
sprite_gubbe_split(12) <= "11111111111111111111001111110010";
sprite_gubbe_split(13) <= "11111111111111111111001111110010";
sprite_gubbe_split(14) <= "11111111111001111111111111110010";
sprite_gubbe_split(15) <= "11111111111001111111111111110010";
sprite_gubbe_split(16) <= "11111111111001111111111111110010";
sprite_gubbe_split(17) <= "11111111111001111111111111110010";
sprite_gubbe_split(18) <= "11111111111001111111111111110010";
sprite_gubbe_split(19) <= "11111001111001111111001111110010";
sprite_gubbe_split(20) <= "11111011111100111111111111110010";
sprite_gubbe_split(21) <= "11111011111100111111111111110010";
sprite_gubbe_split(22) <= "11111111111111111111111111110010";
sprite_gubbe_split(23) <= "11111011111100111111111111110010";
sprite_gubbe_split(24) <= "11100111111110111111111111110010";
sprite_gubbe_split(25) <= "11111111111111111111111111111110";
sprite_gubbe_split(26) <= "11101111111111111111111111110010";
sprite_gubbe_split(27) <= "11111111111111111111111111111110";
sprite_gubbe_split(28) <= "11101111110011111111111111110010";
sprite_gubbe_split(29) <= "11101111111110111111001111110010";
sprite_gubbe_split(30) <= "11111111111111101111001111110010";
sprite_gubbe_split(31) <= "11111111111111111111111111110010";
sprite_gubbe_split(32) <= "11111111111111111111111111111111";
sprite_gubbe_split(33) <= "11110011111100111111111111110010";
sprite_gubbe_split(34) <= "11111110011111111111001111110010";
sprite_gubbe_split(35) <= "11001111101110011111001111110010";
sprite_gubbe_split(36) <= "11001111101110011111001111110010";
sprite_gubbe_split(37) <= "11111111101111111111001111110010";
sprite_gubbe_split(38) <= "11111111111111111111111111110010";
sprite_gubbe_split(39) <= "11111111111111111111111111110010";
sprite_gubbe_split(40) <= "11111111111111111111111111110010";
sprite_gubbe_split(41) <= "11111111111101111111001111110010";
sprite_gubbe_split(42) <= "11111111111101111111001111110010";
sprite_gubbe_split(43) <= "11111111111111111111001111110010";
sprite_gubbe_split(44) <= "11111111111111111111001111110010";
sprite_gubbe_split(45) <= "11111111111111111111001111110010";
sprite_gubbe_split(46) <= "11111111111001111111111111110010";
sprite_gubbe_split(47) <= "11111111111111111111111111111010";
sprite_gubbe_split(48) <= "11111111111001111111111111110010";
sprite_gubbe_split(49) <= "11111111111111111111111111111010";
sprite_gubbe_split(50) <= "11111111111111111111111111111010";
sprite_gubbe_split(51) <= "11111001111111111111111111110010";
sprite_gubbe_split(52) <= "11111011111100111111111111110010";
sprite_gubbe_split(53) <= "11111011111100111111111111110010";
sprite_gubbe_split(54) <= "11111011111100111111111111111110";
sprite_gubbe_split(55) <= "11111011111100111111111111110010";
sprite_gubbe_split(56) <= "11100111111110111111111111110010";
sprite_gubbe_split(57) <= "11101111111100111111001111110010";
sprite_gubbe_split(58) <= "11101111111111111111101111110010";
sprite_gubbe_split(59) <= "11101111110011111111111111110010";
sprite_gubbe_split(60) <= "11101111110011111111111111110010";
sprite_gubbe_split(61) <= "11101111111110111111001111110010";
sprite_gubbe_split(62) <= "11111111111111101111001111110010";
sprite_gubbe_split(63) <= "11111111111111101111001111110010";

process(clk)
variable gubbe: integer :=3;
variable detected: boolean := false;
variable collisionDetected: boolean := false;
begin
	if rising_edge(clk) then
		if rst ='1' then
			x_pos(0) <= 0;
			y_pos(0) <= 200;
			x_pos(1) <= 0;
			y_pos(1) <= 200;
			x_pos(2) <= 0;
			y_pos(2) <= 200;
			x_pos(3) <= 100;
			y_pos(3) <= 200;			
		else		
			if(jump='1') then
				y_pos(gubbe) <= 168;
				sprite_gubbe_aktiv<=sprite_gubbe_jump;
			elsif(duck='1') then
				y_pos(gubbe) <= 232;
				sprite_gubbe_aktiv<=sprite_gubbe_duck;
			else
				y_pos(gubbe) <= 200;
				if split_legs = '1' then
						sprite_gubbe_aktiv<=sprite_gubbe;
				else
						sprite_gubbe_aktiv<=sprite_gubbe_split;
				end if;
			end if;
			
			detected :=false;		
			collisionDetected := false;
			
			if put_box = '1' then
				 if x_pos(0) = 0 then
					x_pos(0) <= 800;
					if next_box ='1' then
						y_pos(0) <= 200;
					else
						y_pos(0) <= 232;
					end if;
				 elsif x_pos(1) = 0 then
					x_pos(1) <= 800;
					if next_box ='1' then
						y_pos(1) <= 200;
					else
						y_pos(1) <= 232;
					end if;
				 elsif x_pos(2) = 0 then
					x_pos(2) <= 800;
					if next_box ='1' then
						y_pos(2) <= 200;
					else
						y_pos(2) <= 232;
					end if;
				 else
				 end if;
			elsif move_box ='1' then
				for i in 2 downto 0 loop
					if x_pos(i)>0 then
						x_pos(i) <= x_pos(i) -1;
					end if;
				end loop;
			end if;

			for i in 2 downto 0 loop
			
				if y>=y_pos(i) and y < (y_pos(i)+spriteSize) then
					if x>= x_pos(i) and x < (x_pos(i)+spriteSize) then
						if sprite_brick( y - y_pos(i) )( x - x_pos(i) ) = '1' then
							spriteVgaRed<="111";				
							spriteVgaGreen<="101";
							spriteVgaBlue<="11";
							detected:= true;
						end if;					
					end if;					
				end if;
						
			end loop;
			
			if y>=y_pos(gubbe) and y < (y_pos(gubbe)+gubbSize) then
				if x>= x_pos(gubbe) and x < (x_pos(gubbe)+spriteSize) then
					if sprite_gubbe_aktiv( y - y_pos(gubbe) )( x - x_pos(gubbe) ) = '1' then
						spriteVgaRed<="111";				
						spriteVgaGreen<="101";
						spriteVgaBlue<="00";
						if detected = true then
							collisionDetected := true;
						end if;
						detected:= true;
					end if;					
				end if;					
			end if;
					
			if detected = true then
				spriteDetected <= '1';
			else
				spriteDetected <= '0';
			end if;
			
			if collisionDetected = true then
				collision <='1';
				else
				collision <='0';
			end if;
		end if;
	end if;
end process;

end Behavioral;

